*KLconst1

*KLayout0

.subckt	bfr1	A	dcin	dcout	q	xin	xout	
B11	4	0	jmod	area=0.5
B21	5	0	jmod	area=0.5
L1	2       4	1.98p    
L2      5	2       1.98p
Ld	DCin 	DCout	7.34p
Lx	Xin	Xout	7.28p
Lin	A	2	2.119p
Lq	2	0	7.511p
Lout	0	q	26.304p

Kx1	Lx	L1	-0.17233
Kx2	Lx	L2	-0.17233
Kxd	Lx	Ld	0.088579
Kd1	Ld	L1	-0.12779
Kd2	Ld	L2	-0.12779
Kind	Lin	Ld	2.638E-4	
Kinx	Lin	Lx	7.711E-5
Kxout	Lx	Lout	-3.194E-5
Kdout	Ld	Lout	-1.522E-5
Kout	Lq	Lout	-0.573
.ends bfr1

.subckt	const1	dcin	dcout	q	xin	xout	
B11	4	0	jmod	area=0.5
B21	5	0	jmod	area=0.5
L1	2       4	2.393p    
L2      5	2       1.885p
Ld	DCin 	DCout	7.369p
Lx	Xin	Xout	7.321p
Lq	2	0	7.412p
Lout	0	q	26.35p

Kx1	Lx	L1	-0.1958
Kx2	Lx	L2	-0.1473 
Kxd	Lx	Ld	0.092378 
Kd1	Ld	L1	-0.1562
Kd2	Ld	L2	-0.0992
Kxout	Lx	Lout	-5.755E-4
Kdout	Ld	Lout	-1.419E-3
Kout	Lq	Lout	-0.57885  
.ends const1

VAC1	AC1	0	SIN(0 811mV 5GHz 100ps 0)
VAC2	0	AC2	SIN(0 811mV 5GHz 150ps 0)
VDC	DC1	0	PWL(0ps 0mv 20ps 1131mV)

Rdc	DC1	d1in	1000 nfree
Rx1	AC1	a1in	1000 nfree
Rx2	AC2	a2in	1000 nfree

Xcon	const1	d1in	dout	q1	a1in	a1out1
X2	bfr1	q1	dout2	dout	out1	a2in	a2out1
X3	bfr1	out1 	dout2	dout3	out2	a1out2	a1out1
X4	bfr1	out2	dout4	dout3	out3	a2out2	a2out1
X5	bfr1	out3	dout4	dout5	out4	a1out2	a1out3
X6	bfr1	out4	dout6	dout5	out5	a2out2	a2out3
X7	bfr1	out5	dout6	dout7	out6	a1out4	a1out3
X8	bfr1	out6	dout8	dout7	out7	a2out4	a2out3
X9	bfr1	out7	dout8	dout9	out8	a1out4	a1out5
X10	bfr1	out8	dout10	dout9	out9	a2out4	a2out5
X11	bfr1	out9	dout10	dout11	out10	0	a1out5
X12	bfr1	out10	0	dout11	0	0	a2out5


.model jmod jj(rtype=1, vg=2.8mV, cap=0.064pF, r0=100, rN=17, icrit=0.1mA, Phi=pi)
.tran 0.2p 3000p 0 0.2p

.print i(Lq|X2)
.print i(Lq|X5)
.print i(Lq|X9)
.print i(Lq|X12)

.end