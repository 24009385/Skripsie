
*JSIM model
**HSTP**
.model jjmod jj(Rtype=1, Vg=2.8mV, Cap=0.064pF, R0=100ohm, Rn=17ohm, Icrit=0.1mA, Phi=pi)
**OPEN**
*.model jjmod jj(Rtype=1, Vg=2.8mV, Cap=0.218pF, R0=200ohm, Rn=17ohm, Icrit=0.1mA)


*** netlist file ***
**** **** **** **** **** **** **** ****+
*** Lib : hstp_komiya_lib
*** Cell: pi_buf3_test
*** View: schematic
*** Jan 16 00:02:30 2022
**** **** **** **** **** **** **** ****

*** pi_buffer3
.subckt pi_buffer3          1          2          3          4          5          6
***         a       din      dout         q       xin      xout
Kxd                Lx         Ld 0.190
Kd2                Ld         L2 -0.133
Kx2                Lx         L2 -0.186
Kx1                Lx         L1 -0.186
Kd1                Ld         L1 -0.133

Bpi2               7         0  jjmod area=0.50
Bpi1               8         0  jjmod area=0.50
Lq1                9        10   0.140pH fcheck
Lq2               10         0   7.780pH fcheck
L2                 7         9   1.590pH fcheck
Lin                1         9   1.230pH fcheck
Lout              10        11  23.420pH fcheck
Lx                 5         6   7.400pH fcheck
Ld                 2         3   7.450pH fcheck
L1                 9         8   1.590pH fcheck
Rout              11         4   1.000pohm nfree
.ends

*** pi_buffer4
.subckt pi_buffer4          1          2          3          4          5          6
***         a       din      dout         q       xin      xout
Kxd                Lx         Ld 0.190
Kd2                Ld         L2 -0.133
Kx2                Lx         L2 -0.186
Kx1                Lx         L1 -0.186
Kd1                Ld         L1 -0.133
Bpi2               7         0  jjmod area=0.50
Bpi1               8         0  jjmod area=0.50
Lq1                9        10   0.140pH fcheck
Lq2               10         0   7.780pH fcheck
L2                 7         9   1.590pH fcheck
Lin                1         9   1.230pH fcheck
Lout              10        11  23.420pH fcheck
Lx                 5         6   7.400pH fcheck
Ld                 2         3   7.450pH fcheck
L1                 9         8   1.590pH fcheck
Rout              11         4   1.000pohm nfree
.ends

*** top cell: pi_buf3_test
Vx2   0    12  SIN(0 811mV 5GHz 150ps 0)
Vdc   13   0   PWL(0ps 0mv 20ps 1131mV)
Vx1   14   0   SIN(0 811mV 5GHz 100ps 0)
Vin   15   0   PWL(0ps 0mV 1ps -5mV 150ps -5mV 350ps -5mV 351ps 5mV 550ps 5mV 551ps -5mV 750ps -5mV 751ps 5mV 950ps 5mV 951ps -5mV 1150ps -5mV 1350ps -5mV 1351ps 5mV 1550ps 5mV 1750ps 5mV )
Rx2               12         8  1000.00ohm nfree
Rdc               13        16  1000.00ohm nfree
Rx1               14        10  1000.00ohm nfree
Rin               15         9  1000.00ohm nfree
XI8        pi_buffer3         17         18          0          0         21          0
*** ("22" "20" "19") mapped to 0
XI5        pi_buffer3         23         24         25         26         27         28
XI6        pi_buffer3         26         24         29         30         21         31
XI7        pi_buffer3         30         18         29         17          0         28
*** ("11") mapped to 0
XI2        pi_buffer3         32         33         34         35          7         36
XI3        pi_buffer3         35         37         34         38         27         39
XI0        pi_buffer3          9         16         40         41         10         36
XI1        pi_buffer3         41         33         40         32          8         39
XI4        pi_buffer4         42         37         25         43          7         31
Lin               38        42   0.000pH fcheck
Lout              43        23   0.000pH fcheck

*** netlist file ***
.tran 0.2ps 3000ps 0ps 0.2ps
.print i(Rx1)
.print i(Rx2)
.print i(Rin)
.print i(Lq2|XI0)
.print i(Lq2|XI1)
.print i(Lq2|XI2)
.print i(Lq2|XI3)
.print i(Lq2|XI4)
.print i(Lq2|XI8)
.print i(Lout)
*** jsim input file ***

*** jsim input file ***