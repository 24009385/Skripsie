
* Example Buffer basic
.subckt	bfr1	A	dcin	dcout	q	xin	xout	

B11	4	0	jmod	area=0.5
B21	5	0	jmod	area=0.5
L1	2       4	1.59p    
L2      5	2       1.59p
Ld	DCin 	DCout	6.8p
Lx	Xin	Xout	6.7p
Lin	A	2	1.22p
Lq	2	0	7.93p
Lout	q	0	31p

Kx1	Lx	L1	-0.186
Kx2	Lx	L2	-0.186
Kxd	Lx	Ld	0.190
Kd1	Ld	L1	-0.133
Kd2	Ld	L2	-0.133
Kind	Lin	Ld	5.063E-4	
Kinx	Lin	Lx	3.145E-5
Kxout	Lx	Lout	2.02E-3
Kdout	Ld	Lout	2.69E-5
Kout	Lq	Lout	0.691
.ends bfr1

VAC1	AC1	0	SIN(0 811mV 5GHz 100ps 0)
VAC2	0	AC2	SIN(0 811mV 5GHz 150ps 0)
VDC	DC1	0	PWL(0ps 0mv 20ps 1131mV)
Vin	In1	0	PWL(0ps 0mV 1ps -5mV 150ps -5mV 350ps -5mV 351ps 5mV 550ps 5mV 551ps -5mV 750ps -5mV 751ps 5mV 950ps 5mV 951ps -5mV 1150ps -5mV 1350ps -5mV 1351ps 5mV 1550ps 5mV 1750ps 5mV )

Rin	In1	1	1000 nfree
Rdc	DC1	d1in	1000 nfree
Rx1	AC1	a1in	1000 nfree	
Rx2	AC2	a2in	1000 nfree

*X	name	a	dcin	dcout	q	xin	xout

Xbfr1  	bfr1	1	d1in	d1out	bfr1out	a1in	a1out	
Xbfr2   bfr1	bfr1out	d2in	d1out	bfr2out	a2in	a2out	
Xbfr3 	bfr1	bfr2out	d2in	d2out	bfr3out	0	a1out	
Xbfr4	bfr1	bfr3out	0	d2out	Out	0	a2out	

Lyout	Out	0	0 



.model jmod jj(rtype=1, vg=2.8mV, cap=0.064pF, r0=100, rN=17, icrit=0.1mA, Phi=pi)
.tran 0.2p 3000p 0 0.2p
.print I(Lq|Xbfr1)
.print I(Lq|Xbfr2)
.print I(Lq|Xbfr3)
.print I(Lq|Xbfr4)
.print i(Lout|Xbfr1)
.print i(Rx1)
.print i(Rx2)
.print i(Rin)
.print i(Lyout)
.end