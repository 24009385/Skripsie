* OR3

.subckt	bias	DCin	DCout	Xin	Xout
Lb0	DCin 	DCout	6p
Lb1	Xin	Xout	6p
.ends bias

.subckt OR3	DCin	DCout	InA	InB	InC	q	Xin	Xout
Xb1	bias	DCin	dout1	Xin	a1out1
Xbfr1	bfr1	InA	dout1	dout2	q1	a1out1	a1out2
Xconst1	const1	dout2	dout3	q4	a1out2	a1out3
Xbfr2	bfr1	InB	dout3	dout4	q2	a1out3	a1out4
Xconst2	const1	dout4	dout5	q5	a1out4	a1out5
Xbfr3	bfr1	InC	dout5	dout6	q3	a1out5	a1out6
Xb2	bias	dout6	DCout	a1out6	Xout

La	q1	qm	16p
Lb	q2	qm	16p
Lc	q3	qm	16p
Ld	q4	qm	16p
Le	q5	qm	16p
Lo	qm	q	0.17p
.ends OR3

.subckt	const1	dcin	dcout	q	xin	xout	
.model jmod jj(rtype=1, vg=2.8mV, cap=0.064pF, r0=100, rN=17, icrit=0.1mA, Phi=pi)
B11	4	0	jmod	area=0.5
B21	5	0	jmod	area=0.5
L1	2       4	1.6p    
L2      5	2       1.75p
Ld	DCin 	DCout	6.6p
Lx	Xin	Xout	6.6p
Lq	2	0	8.2p
Lout	q	0	30.5p
Kx1	Lx	L1	-0.22
Kx2	Lx	L2	-0.26
Kxd	Lx	Ld	0.290
Kd1	Ld	L1	-0.168
Kd2	Ld	L2	-0.208
Kxout	Lx	Lout	-2.42E-4
Kdout	Ld	Lout	-5.49E-4
Kout	Lq	Lout	-0.8
.ends const1


.subckt	bfr1	A	dcin	dcout	q	xin	xout	
B11	4	0	jmod	area=0.5
B21	5	0	jmod	area=0.5
L1	2       4	1.59p    
L2      5	2       1.59p
Ld	DCin 	DCout	6.8p
Lx	Xin	Xout	6.7p
Lin	A	2	1.22p
Lq	2	0	7.93p
Lout	0	q	31p
Kx1	Lx	L1	-0.186
Kx2	Lx	L2	-0.186
Kxd	Lx	Ld	0.190
Kd1	Ld	L1	-0.133
Kd2	Ld	L2	-0.133
Kind	Lin	Ld	5.063E-4	
Kinx	Lin	Lx	3.145E-5
Kxout	Lx	Lout	2.02E-3
Kdout	Ld	Lout	2.69E-5
Kout	Lq	Lout	-0.691
.ends bfr1


VAC1	AC1	0	SIN(0 811mV 5GHz 100ps 0)
VAC2	0	AC2	SIN(0 811mV 5GHz 150ps 0)
VDC	DC1	0	PWL(0ps 0mv 20ps 1131mV)

VinA	InA	0	PWL(0ps 0mV 1ps -5mV 	150ps -5mV 350ps -5mV 	351ps -5mV 550ps -5mV		551ps -5mV 750ps -5mV 		751ps -5mV 950ps -5mV 							951ps 5mV 1150ps 5mV 	1151ps 5mv 1350ps 5mV 		1351ps 5mV 1550ps 5mV 		1151ps 5mV 1750ps 5mV	1751ps -5mV)
*Above (00001111)

VinB	InB	0	PWL(0ps 0mV 1ps -5mV 	150ps -5mV 350ps -5mV 	351ps -5mV 550ps -5mV		551ps 5mV 750ps 5mV 		751ps 5mV 950ps 5mV 							951ps -5mV 1150ps -5mV 	1151ps -5mv 1350ps -5mV 	1351ps 5mV 1550ps 5mV 		1151ps 5mV 1750ps 5mV		1751ps -5mV)
*Above (00110011)

VinC	InC	0	PWL(0ps 0mV 1ps -5mV 	150ps -5mV 350ps -5mV 	351ps 5mV 550ps 5mV		551ps -5mV 750ps -5mV 		751ps 5mV 950ps 5mV 							951ps -5mV 1150ps -5mV 	1151ps 5mv 1350ps 5mV 		1351ps -5mV 1550ps -5mV 	1151ps 5mV 1750ps 5mV		1751ps -5mV)
*Above (01010101)


RinA	InA	A	1000 nfree
RinB	InB  	B	1000 nfree
RinC	InC	C	1000 nfree

Rdc	DC1	d1in	1000 nfree
Rx1	AC1	a1in	1000 nfree
Rx2	AC2	a2in	1000 nfree

XA	bfr1	A	d1in	dout1	ao	a1in	a1out1
XB	bfr1	B	dout1	dout2	bo	a1out1	a1out2
XC	bfr1	C	dout2	dout3	co	a1out2	a1out3

XAND	OR3	dout4	dout3	ao	bo	co	q0	a2in	a2out1

X1	bfr1	q0	dout4	dout5	q1	0	a1out3

X2	bfr1	q1	0	dout5	0	0	a2out1

.model jmod jj(rtype=1, vg=2.8mV, cap=0.064pF, r0=100, rN=17, icrit=0.1mA, Phi=pi)
.tran 0.2p 3000p 0 0.2p

.print i(RinA)
.print i(RinB)
.print i(RinC)

.print i(Lq|X1)
.print i(Lq|X2)
.end