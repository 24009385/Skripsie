*FAt2

.subckt	bias 	DCin	DCout	Xin	Xout
Lb0	DCin 	DCout	0
Lb1	Xin	Xout	0
.ends bias

.subckt OR2	DCin	DCout	InA	InB	q	Xin	Xout
Xbfr1	bfr1	InA	DCin	d1out	q1	Xin	a1out	
Xconst	const1	d1out	d2out	q2	a1out	a2out
Xbfr3	bfr1	InB	d2out	DCout	q3	a2out	Xout
La	q1	q	16p
Lb	q2	q	16p
Lc	q3	q	16p
.ends OR2

.subckt OR3	DCin	DCout	InA	InB	InC	q	Xin	Xout
Xb1	bias	DCin	dout1	Xin	a1out1
Xbfr1	bfr1	InA	dout1	dout2	q1	a1out1	a1out2
Xconst1	const1	dout2	dout3	q4	a1out2	a1out3
Xbfr2	bfr1	InB	dout3	dout4	q2	a1out3	a1out4
Xconst2	const1	dout4	dout5	q5	a1out4	a1out5
Xbfr3	bfr1	InC	dout5	dout6	q3	a1out5	a1out6
Xb2	bias	dout6	DCout	a1out6	Xout

La	q1	qm	16p
Lb	q2	qm	16p
Lc	q3	qm	16p
Ld	q4	qm	16p
Le	q5	qm	16p
Lo	qm	q	0.17p
.ends OR3

.subckt	const1	dcin	dcout	q	xin	xout	
.model jmod jj(rtype=1, vg=2.8mV, cap=0.064pF, r0=100, rN=17, icrit=0.1mA, Phi=pi)
B11	4	0	jmod	area=0.5
B21	5	0	jmod	area=0.5
L1	2       4	1.6p    
L2      5	2       1.75p
Ld	DCin 	DCout	6.6p
Lx	Xin	Xout	6.6p
Lq	2	0	8.2p
Lout	q	0	30.5p

Kx1	Lx	L1	-0.22
Kx2	Lx	L2	-0.26
Kxd	Lx	Ld	0.290
Kd1	Ld	L1	-0.168
Kd2	Ld	L2	-0.208
Kxout	Lx	Lout	-2.42E-4
Kdout	Ld	Lout	-5.49E-4
Kout	Lq	Lout	-0.6
.ends const1

.subckt	const0	dcin	dcout	q	xin	xout	
B11	4	0	jmod	area=0.5
B21	5	0	jmod	area=0.5
L1	2       4	1.6p    
L2      5	2       1.75p
Ld	DCin 	DCout	6.6p
Lx	Xin	Xout	6.6p
Lq	2	0	8.2p
Lout	q	0	30.5p
Kx1	Lx	L1	-0.22
Kx2	Lx	L2	-0.26
Kxd	Lx	Ld	0.290
Kd1	Ld	L1	-0.168
Kd2	Ld	L2	-0.208
Kxout	Lx	Lout	-2.42E-4
Kdout	Ld	Lout	-5.49E-4
Kout	Lq	Lout	0.6
.ends const0

.subckt AND2	DCin	DCout	InA	InB	q	Xin	Xout
Xbfr1  	bfr1	InA	DCin	d1out	q1	Xin	a1out
Xconst	const0	d1out 	d2out	q2	a1out	a2out
Xbfr3  	bfr1	InB	d2out	DCout	q3	a2out	Xout
La	q1	q	10p
Lb	q2	q	60p
Lc	q3	q	10p
.ends AND2

.subckt AND3	DCin	DCout	InA	InB	InC	q	Xin	Xout
Xb1	bias	DCin	dout1	Xin	a1out1
Xbfr1	bfr1	InA	dout1	dout2	q1	a1out1	a1out2
Xconst1	const0	dout2	dout3	q4	a1out2	a1out3
Xbfr2	bfr1	InB	dout3	dout4	q2	a1out3	a1out4
Xconst2	const0	dout4	dout5	q5	a1out4	a1out5
Xbfr3	bfr1	InC	dout5	dout6	q3	a1out5	a1out6
Xb2	bias	dout6	DCout	a1out6	Xout

La	q1	qm	16p
Lb	q2	qm	16p
Lc	q3	qm	16p
Ld	q4	qm	16p
Le	q5	qm	16p
Lo	qm	q	0.17p
.ends AND3

.subckt	splitWB	A	dcin	dcout	q	xin	xout	
B11	4	0	jmod	area=0.5
B21	5	0	jmod	area=0.5
L1	2       4	1.59p    
L2      5	2       1.59p
Ld	8 	9	6.8p
Lx	10	11	6.7p
Lin	A	2	1.22p
Lq	2	0	7.93p
Lout	q	0	31p
Lb1	9	DCout 	0
Lb0	DCin 	8	0
Lb3	11	Xout 	0p
Lb2	Xin 	10	0p
Kx1	Lx	L1	-0.186
Kx2	Lx	L2	-0.186
Kxd	Lx	Ld	0.190
Kd1	Ld	L1	-0.133
Kd2	Ld	L2	-0.133
Kind	Lin	Ld	5.063E-4	
Kinx	Lin	Lx	3.145E-5
Kxout	Lx	Lout	2.02E-3
Kdout	Ld	Lout	2.69E-5
Kout	Lq	Lout	0.691
.ends splitWB

.subckt branch	a	b	q
Lq	1	q	0.17p
Lb	b	1	10.4p
La	a	1	10.4p
.ends branch

.subckt split	A	DCin	DCout	q0	q1	Xin	Xout
Xsplit 	splitWB	A	DCin	DCout	out	Xin	Xout
Xq	branch	q0 	q1	out
.ends split

.subckt	bfr1	A	dcin	dcout	q	xin	xout	
B11	4	0	jmod	area=0.5
B21	5	0	jmod	area=0.5
L1	2       4	1.59p    
L2      5	2       1.59p
Ld	DCin 	DCout	6.8p
Lx	Xin	Xout	6.7p
Lin	A	2	1.22p
Lq	2	0	7.93p
Lout	0	q	31p
Kx1	Lx	L1	-0.186
Kx2	Lx	L2	-0.186
Kxd	Lx	Ld	0.190
Kd1	Ld	L1	-0.133
Kd2	Ld	L2	-0.133
Kind	Lin	Ld	5.063E-4	
Kinx	Lin	Lx	3.145E-5
Kxout	Lx	Lout	2.02E-3
Kdout	Ld	Lout	2.69E-5
Kout	Lq	Lout	-0.691
.ends bfr1

.subckt	bfrN	A	dcin	dcout	q	xin	xout
B11	4	0	jmod	area=0.5
B21	5	0	jmod	area=0.5
L1	2       4	1.59p    
L2      5	2       1.59p
Ld	DCin 	DCout	6.8p
Lx	Xin	Xout	6.7p
Lin	A	2	1.22p
Lq	2	0	7.93p
Lout	0	q	31p
Kx1	Lx	L1	-0.186
Kx2	Lx	L2	-0.186
Kxd	Lx	Ld	0.190
Kd1	Ld	L1	-0.133
Kd2	Ld	L2	-0.133
Kind	Lin	Ld	5.063E-4	
Kinx	Lin	Lx	3.145E-5
Kxout	Lx	Lout	2.02E-3
Kdout	Ld	Lout	2.69E-5
Kout	Lq	Lout	0.691
.ends bfrN

VAC1	AC1	0	SIN(0 811mV 5GHz 100ps 0)
VAC2	0	AC2	SIN(0 811mV 5GHz 150ps 0)
VDC	DC1	0	PWL(0ps 0mv 20ps 1131mV)

VinA	InA	0	PWL(0ps 0mV 1ps -5mV 	150ps -5mV 350ps -5mV 	351ps -5mV 550ps -5mV		551ps -5mV 750ps -5mV 		751ps -5mV 950ps -5mV 							951ps 5mV 1150ps 5mV 	1151ps 5mv 1350ps 5mV 		1351ps 5mV 1550ps 5mV 		1151ps 5mV 1750ps 5mV	1751ps -5mV)
*Above (00001111)

VinB	InB	0	PWL(0ps 0mV 1ps -5mV 	150ps -5mV 350ps -5mV 	351ps -5mV 550ps -5mV		551ps 5mV 750ps 5mV 		751ps 5mV 950ps 5mV 							951ps -5mV 1150ps -5mV 	1151ps -5mv 1350ps -5mV 	1351ps 5mV 1550ps 5mV 		1151ps 5mV 1750ps 5mV		1751ps -5mV)
*Above (00110011)

VinC	InC	0	PWL(0ps 0mV 1ps -5mV 	150ps -5mV 350ps -5mV 	351ps 5mV 550ps 5mV		551ps -5mV 750ps -5mV 		751ps 5mV 950ps 5mV 							951ps -5mV 1150ps -5mV 	1151ps 5mv 1350ps 5mV 		1351ps -5mV 1550ps -5mV 	1151ps 5mV 1750ps 5mV		1751ps -5mV)
*Above (01010101)

RinA	InA	A	1000 nfree
RinB	InB  	B	1000 nfree
RinC	InC	C	1000 nfree

Rdc	DC1	d1in	1000 nfree
Rx1	AC1	a1in	1000 nfree
Rx2	AC2	a2in	1000 nfree


*XsplitA	split	In1	DCin	d1out	q01	q11	Xin1	a1out1
XsA	split	A	d1in	dout1	qa0	qa1	a1in	a1out1
XsB	split	B	dout1	dout2	qb0	qb1	a1out1	a1out2
XsC	split	C	dout2	dout3	qc0	qc1	a1out2	a1out3

XA1	bfr1	qa0	dout9	dout8	qa2	a2out5	a2out6
XA2	bfr1	qa1	dout8	dout7	qa3	a2out4	a2out5
XB1	bfr1	qb0	dout7	dout6	qb2	a2out3	a2out4
XB2	bfr1	qb1	dout6	dout5	qb3	a2out2	a2out3
XC1	bfr1	qc0	dout5	dout4	qc2	a2out1	a2out2
XC2	bfr1	qc1	dout4	dout3	qc3	a2in	a2out1

XsA1	split	qa2	dout9	dout10	qa4	qa5	a1out4	a1out3
XsA2	split	qa3	dout10	dout11	qa6	qa7	a1out5	a1out4
XsB1	split	qb2	dout11	dout12	qb4	qb5	a1out6	a1out5
XsB2	split	qb3	dout12	dout13	qb6	qb7	a1out7	a1out6
XsC1	split	qc2	dout13	dout14	qc4	qc5	a1out8	a1out7
XsC2	bfr1	qc3	dout14	dout15	qc6	a1out9	a1out8

XssA1	bfr1	qa4	dout16	dout15	qao1	a2out7	a2out6
XssA2	bfr1	qa5	dout17	dout16	qao2	a2out8	a2out7
XssA3	bfr1	qa6	dout18	dout17	qao3	a2out9	a2out8
XssA4	bfr1	qa7	dout19	dout18	qao4	a2out10	a2out9
XssB1	bfr1	qb4	dout20	dout19	qbo1	a2out11	a2out10
XssB2	bfr1	qb5	dout21	dout20	qbo2	a2out12	a2out11
XssB3	bfr1	qb6	dout22	dout21	qbo3	a2out13	a2out12
XssB4	bfr1	qb7	dout23	dout22	qbo4	a2out14	a2out13
XssC1	bfr1	qc4	dout24	dout23	qco1	a2out15	a2out14
XssC2	bfr1	qc5	dout25	dout24	qco2	a2out16	a2out15
XssC3	bfr1	qc6	dout26	dout25	qco3	a2out17	a2out16

Xor1	OR2	dout32	dout33	qao1	qbo1	oi1	a1out9	a1out10
Xand1	AND2	dout31	dout32	qao2	qbo2	oi2	a1out10	a1out11
Xbfr1	bfr1	qco3	dout30	dout31	oi3	a1out11	a1out12

Xo31	OR2	dout29	dout30	qao3	qbo3	oi4	a1out12	a1out13
Xob1	bfr1	qco1	dout28	dout29	oi5	a1out13	a1out14

Xa31	AND2	dout27	dout28	qao4	qbo4	oi6	a1out14	a1out15
Xab1	bfr1	qco2	dout26	dout27	oi7	a1out15	a1out16

Xaz1	bfr1	oi1	dout34	dout33	o1	a2out17	a2out18		
Xaz2	bfr1	oi2	dout35	dout34	o2	a2out18	a2out19		
Xaz3	bfr1	oi3	dout36	dout35	o3	a2out19 a2out20
Xaz4	bfr1	oi4	dout37	dout36	o4	a2out20	a2out21	
Xaz5	bfr1	oi5	dout38	dout37	o5	a2out21	a2out22
Xaz6	bfr1	oi6	dout39	dout38	o6	a2out22	a2out23
Xaz7	bfr1	oi7	dout40	dout39	o7	a2out23	a2out24

Xo32	OR2	dout40	dout41	o4	o5	op1	a1out17	a1out16
Xa32	AND2	dout41	dout42	o6	o7	op2	a1out18	a1out17
Xand2	AND2	dout42	dout43	o1	o3	op3	a1out19	a1out18
Xbfr3	bfr1	o2	dout43	dout44	op4	a1out20	a1out19


Xe1	bfr1	op1	dout45	dout44	o11	a2out25	a2out24
Xe2	bfr1	op2	dout46	dout45	o21	a2out26	a2out25
Xe3	bfr1	op3	dout47	dout46	o31	a2out27	a2out26
Xe4	bfr1	op4	dout48	dout47	o41	a2out28	a2out27

Xor3	OR2	dout48	dout49	o31	o41	o14	a1out20	a1out21
Xh1	bfr1	o21	dout49	dout50	o34	a1out21	a1out22
Xh2	bfr1	o11	dout50	dout51	o24	a1out22	a1out23


*Done until here


Xi1	bfr1	o14	dout52	dout51	o15	a2out28	a2out29	
Xi2	bfr1	o24	dout53	dout52	o25	a2out29	a2out30	
Xi3	bfr1	o34	dout54	dout53	o35	a2out30	a2out31	

Xj1	bfrN	o15	dout54	dout55	o16	a1out24	a1out23
Xj2	bfr1	o25	dout55	dout56	o26	a1out25	a1out24	
Xj3	bfr1	o35	dout56	dout57	o36	a1out26	a1out25	

Xisplt	split	o16	dout58	dout57	o171	o172	a2out32	a2out31
Xis1	bfr1	o26	dout59	dout58	o27	a2out33	a2out32
Xis2	bfr1	o36	dout60	dout59	o37	a2out34	a2out33

Xk1	bfrN	o171	dout60	dout61	o181	a1out26	a1out27	
Xk2	bfr1	o172	dout61	dout62	o182	a1out27	a1out28	
Xk3	bfr1	o27	dout62	dout63	o28	a1out28	a1out29	
Xk4	bfr1	o37	dout63	dout64	o38	a1out29	a1out30	

XL1	bfr1	o181	dout65	dout64	o191	a2out34	a2out35
XL2	bfr1	o182	dout66	dout65	o192	a2out35	a2out36	
XL3	bfr1	o28	dout67	dout66	o29	a2out36	a2out37	
XL4	bfr1	o38	dout68	dout67	o39	a2out37	a2out38	

Xm1	bfr1	o191	dout68	dout69	o110	a1out31	a1out30
*Xm1 is the Cout
Xand4	AND2	dout69	dout70	o192	o29	o210	a1out32	a1out31
Xm2	bfr1	o39	dout70	dout71	o310	a1out33	a1out32

Xn1	bfr1	o110	dout72	dout71	Cout1	a2out39	a2out38
Xn2	bfr1	o210	dout73	dout72	out1	a2out40	a2out39
Xn3	bfr1	o310	dout74	dout73	out2	a2out41	a2out40

XCout1	bfr1	Cout1	dout74	dout75	Cout2	a1out33	a1out34
Xor4	OR2	dout75	dout76	out1	out2	Sout1	a1out34	0

Xcout	bfr1	Cout2	dout77	dout76	Cout	a2out41	a2out42
Xsum	bfr1	Sout1	0	dout77	Sout	a2out42	0

.model jmod jj(rtype=1, vg=2.8mV, cap=0.064pF, r0=100, rN=17, icrit=0.1mA, Phi=pi)
.tran 0.2p 3000p 0 0.2p

.print i(Lq|Xcout)
.print i(lq|Xsum)

.end