* AND3

.subckt	bias	DCin	DCout	Xin	Xout
Lb0	DCin 	DCout	6p
Lb1	Xin	Xout	6p
.ends bias

.subckt AND3	DCin	DCout	InA	InB	InC	q	Xin	Xout
Xb1	bias	DCin	dout1	Xin	a1out1
Xbfr1	bfr1	InA	dout1	dout2	q1	a1out1	a1out2
Xconst1	const0	dout2	dout3	q4	a1out2	a1out3
Xbfr2	bfr1	InB	dout3	dout4	q2	a1out3	a1out4
Xconst2	const0	dout4	dout5	q5	a1out4	a1out5
Xbfr3	bfr1	InC	dout5	dout6	q3	a1out5	a1out6
Xb2	bias	dout6	DCout	a1out6	Xout

La	q1	qm	16p
Lb	q2	qm	16p
Lc	q3	qm	16p
Ld	q4	qm	16p
Le	q5	qm	16p
Lo	qm	q	0.17p
.ends AND3

.subckt	const0	dcin	dcout	q	xin	xout	
B11	4	0	jmod	area=0.5
B21	5	0	jmod	area=0.5
L1	2       4	1.877p    
L2      5	2       2.402p
Ld	DCin 	DCout	7.369p
Lx	Xin	Xout	7.321p
Lq	2	0	7.412p
Lout	0	q	26.35p

Kx1	Lx	L1	-0.14702 
Kx2	Lx	L2	-0.196 
Kxd	Lx	Ld	0.092378 
Kd1	Ld	L1	-0.098079 
Kd2	Ld	L2	-0.15714
Kxout	Lx	Lout	-5.620E-4
Kdout	Ld	Lout	-1.441E-3
Kout	Lq	Lout	-0.57885  
.ends const0

.subckt	bfr1	A	dcin	dcout	q	xin	xout	
B11	4	0	jmod	area=0.5
B21	5	0	jmod	area=0.5
L1	2       4	1.98p    
L2      5	2       1.98p
Ld	DCin 	DCout	7.34p
Lx	Xin	Xout	7.28p
Lin	A	2	2.119p
Lq	2	0	7.511p
Lout	0	q	26.304p

Kx1	Lx	L1	-0.17233
Kx2	Lx	L2	-0.17233
Kxd	Lx	Ld	0.088579
Kd1	Ld	L1	-0.12779
Kd2	Ld	L2	-0.12779
Kind	Lin	Ld	2.638E-4	
Kinx	Lin	Lx	7.711E-5
Kxout	Lx	Lout	-3.194E-5
Kdout	Ld	Lout	-1.522E-5
Kout	Lq	Lout	-0.573
.ends bfr1


VAC1	AC1	0	SIN(0 811mV 5GHz 100ps 0)
VAC2	0	AC2	SIN(0 811mV 5GHz 150ps 0)
VDC	DC1	0	PWL(0ps 0mv 20ps 1131mV)

VinA	InA	0	PWL(0ps 0mV 1ps -5mV 	150ps -5mV 350ps -5mV 	351ps -5mV 550ps -5mV		551ps -5mV 750ps -5mV 		751ps -5mV 950ps -5mV 							951ps 5mV 1150ps 5mV 	1151ps 5mv 1350ps 5mV 		1351ps 5mV 1550ps 5mV 		1151ps 5mV 1750ps 5mV	1751ps -5mV)
*Above (00001111)

VinB	InB	0	PWL(0ps 0mV 1ps -5mV 	150ps -5mV 350ps -5mV 	351ps -5mV 550ps -5mV		551ps 5mV 750ps 5mV 		751ps 5mV 950ps 5mV 							951ps -5mV 1150ps -5mV 	1151ps -5mv 1350ps -5mV 	1351ps 5mV 1550ps 5mV 		1151ps 5mV 1750ps 5mV		1751ps -5mV)
*Above (00110011)

VinC	InC	0	PWL(0ps 0mV 1ps -5mV 	150ps -5mV 350ps -5mV 	351ps 5mV 550ps 5mV		551ps -5mV 750ps -5mV 		751ps 5mV 950ps 5mV 							951ps -5mV 1150ps -5mV 	1151ps 5mv 1350ps 5mV 		1351ps -5mV 1550ps -5mV 	1151ps 5mV 1750ps 5mV		1751ps -5mV)
*Above (01010101


RinA	InA	A	1000 nfree
RinB	InB  	B	1000 nfree
RinC	InC	C	1000 nfree

Rdc	DC1	d1in	1000 nfree
Rx1	AC1	a1in	1000 nfree
Rx2	AC2	a2in	1000 nfree


XA1	bfr1	A	d1in	dout1	ao	a1in	a1out1
XB1	bfr1	B	dout1	dout2	bo	a1out1	a1out2
XC1	bfr1	C	dout2	dout3	co	a1out2	a1out3

XA2	bfr1	ao	dout4	dout3	ao1	a2in	a2out1
XB2	bfr1	bo	dout5	dout4	bo1	a2out1	a2out2
XC2	bfr1	co	dout6	dout5	co1	a2out2	a2out3

XA3	bfr1	ao1	dout6	dout7	ao2	a1out4	a1out3	
XB3	bfr1	bo1	dout7	dout8	bo2	a1out5	a1out4
XC3	bfr1	co1	dout8	dout9	co2	a1out6	a1out5

XA4	bfr1	ao2	dout10	dout9	ao3	a2out4	a2out3
XB4	bfr1	bo2	dout11	dout10	bo3	a2out5	a2out4
XC4	bfr1	co2	dout12	dout11	co3	a2out6	a2out5

XAND1	AND3	dout12	dout13	ao3	bo3	co3	qa	a1out6	a1out7

X1	bfr1	qa	dout14	dout13	out	a2out6	0
X2	bfr1	out	dout14	0	0	0	a1out7


.model jmod jj(rtype=1, vg=2.8mV, cap=0.064pF, r0=100, rN=17, icrit=0.1mA, Phi=pi)
.tran 0.2p 3000p 0 0.2p


.print i(Lq|X1)
.print i(Lq|X2)

.end