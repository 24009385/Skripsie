* Boost1

.subckt	bfr1	A	dcin	dcout	q	xin	xout	
.model jmod jj(rtype=1, vg=2.8mV, cap=0.064pF, r0=100, rN=17, icrit=0.1mA, Phi=pi)
B11	4	0	jmod	area=0.5
B21	5	0	jmod	area=0.5
L1	2       4	1.59p    
L2      5	2       1.59p
Ld	DCin 	DCout	6.8p
Lx	Xin	Xout	6.7p
Lin	A	2	1.22p
Lq	2	0	7.93p
Lout	q	0	30p

Kx1	Lx	L1	-0.186
Kx2	Lx	L2	-0.186
Kxd	Lx	Ld	0.190
Kd1	Ld	L1	-0.133
Kd2	Ld	L2	-0.133
Kind	Lin	Ld	5.063E-4	
Kinx	Lin	Lx	3.145E-5
Kxout	Lx	Lout	2.02E-3
Kdout	Ld	Lout	2.69E-5
Kout	Lq	Lout	0.691
.ends bfr1

.subckt	boost	A	dcin	dcout	q	xin	xout	
.model jmod jj(rtype=1, vg=2.8mV, cap=0.064pF, r0=100, rN=17, icrit=0.1mA, Phi=pi)
Lin	A	1	0.17p

Lina	1	2	4.9p
L11	2       4	1.45p    
L12     6	2	1.41p
B11	4	0	jmod	area=0.5
B12	6	0	jmod	area=0.5
Lqa	2	0	8.44p

Linb	1	3	4.9p
L21	3       5	1.45p    
L22     7	3	1.41p
B21	5	0	jmod	area=0.5
B22	7	0	jmod	area=0.5
Lqb	3	0	8.44p

Ld	DCin 	DCout	13.11p
Lx	Xin	Xout	12.97p

Lout	0	q	63.8p

Kxa1	Lx	L11	-0.182
Kxa2	Lx	L12	-0.181
Kxb1	Lx	L21	-0.181
Kxb2	Lx	L22	-0.181

Kxd	Lx	Ld	0.287

Kda1	Ld	L11	-0.141
Kda2	Ld	L12	-0.1417
Kdb1	Ld	L21	-0.141
Kdb2	Ld	L22	-0.1408

KoutA	Lout	Lqa	0.428
KoutB	Lout	Lqb	0.38

Kdqa	Ld 	Lqa	-1.55E-3
Kxqa	Lx	Lqa	-1.265E-3
Kdqb	Ld	Lqb	1.873E-3
Kxqb	Lx	Lqb	1.546E-3

Kxout	Lx	Lout	7.708E-4
Kdout	Ld	Lout	1.12E-3

Kdina	Ld	Lina	-5.063E-3	
Kdinb	Ld	Linb	5.863E-3
Kxina	Lx	Lina	-8.845E-3
Kxinb	Lx	Linb	8.745E-3
.ends boost


VAC1	AC1	0	SIN(0 811mV 5GHz 100ps 0)
VAC2	0	AC2	SIN(0 811mV 5GHz 150ps 0)
VDC	DC1	0	PWL(0ps 0mv 20ps 1131mV)

Vin1	In1	0	PWL(0ps 0mV 1ps -5mV 150ps -5mV 350ps -5mV 351ps 5mV 550ps 5mV 551ps -5mV 750ps -5mV 751ps 5mV 950ps 5mV 951ps -5mV 1150ps -5mV 1350ps -5mV 1351ps 5mV 1550ps 5mV 1750ps 5mV )

Rin1	In1	1	1000 nfree
Rdc	DC1	d1in	1000 nfree
Rx1	AC1	a1in	1000 nfree
Rx2	AC2	a2in	1000 nfree

X1  	bfr1	1	d1in	d1out	q0	a1in	0
Ljoin	q0	0	0
X2  	boost	q1	0	d1out	out	a2in	0

Lout 	out	0	0

.tran 0.25p 3000p 0 0.25p
.print i(Lq|X1)
.print i(Lout)
.print i(Ljoin)
.print i(Lqb|X2)
.print i(Lqa|X2)
.print i(Lin|X2)
.print i(Lina|X2)
.print i(Linb|X2)
.end

