
*bfr2

.subckt	bfr2	A	dcin	dcout	q0	q1	xin	xout
B11	4	0	jmod	area=0.5
B21	5	0	jmod	area=0.5
L1	2       4	1.59p    
L2      5	2       1.59p
Ld	DCin 	DCout	6.8p
Lx	Xin	Xout	6.7p
Lin	A	2	1.22p
Lq	2	0	7.93p
Lout	0	1	30p
Lj	1	9	0.8p
Lo1	9	q0	14p
Lo2	9	q1	14p


Kx1	Lx	L1	-0.23
Kx2	Lx	L2	-0.23
Kxd	Lx	Ld	0.2322
Kd1	Ld	L1	-0.16
Kd2	Ld	L2	-0.16
Kind	Lin	Ld	5.063E-4	
Kinx	Lin	Lx	3.145E-5
Kxout	Lx	Lout	2.02E-3
Kdout	Ld	Lout	2.69E-5
Kout	Lq	Lout	-0.691
.ends bfr2

VAC1	AC1	0	SIN(0 811mV 5GHz 100ps 0)
VDC	DC1	0	PWL(0ps 0mv 20ps 1131mV)

Vin	In1	0	PWL(0ps 0mV 1ps -5mV 150ps -5mV 350ps -5mV 351ps 5mV 550ps 5mV 551ps -5mV 750ps -5mV 751ps 5mV 950ps 5mV 951ps -5mV 1150ps -5mV 1350ps -5mV 1351ps 5mV 1550ps 5mV 1750ps 5mV )

Rin	In1	1	1000	0
Rdc	DC1	d1in	1000	0	
Rx1	AC1	a1in	1000	0


Xbfr1	bfr2	1	d1in	0	o1	o2	a1in	0

Lout1	o1	0	0	
Lout2	o2	0	0



.model jmod jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rN=16, icrit=0.1mA)
.tran 0.25p 4000p 0 0.25p
.print i(Lout1)
.print i(Lout2)
.print i(Rin)
.end