* Split Circuit 

.subckt	splitWB	A	dcin	dcout	q	xin	xout	
B11	4	0	jmod	area=0.5
B21	5	0	jmod	area=0.5
L1	2       4	1.59p    
L2      5	2       1.59p
Ld	8 	9	6.8p
Lx	10	11	6.7p
Lin	A	2	1.22p
Lq	2	0	7.93p
Lout	q	0	31p
Lb1	9	DCout 	0
Lb0	DCin 	8	0
Lb3	11	Xout 	0p
Lb2	Xin 	10	0p
Kx1	Lx	L1	-0.186
Kx2	Lx	L2	-0.186
Kxd	Lx	Ld	0.190
Kd1	Ld	L1	-0.133
Kd2	Ld	L2	-0.133
Kind	Lin	Ld	5.063E-4	
Kinx	Lin	Lx	3.145E-5
Kxout	Lx	Lout	2.02E-3
Kdout	Ld	Lout	2.69E-5
Kout	Lq	Lout	0.691
.ends splitWB

.subckt	bfr1	A	dcin	dcout	q	xin	xout	
B11	4	0	jmod	area=0.5
B21	5	0	jmod	area=0.5
L1	2       4	1.59p    
L2      5	2       1.59p
Ld	DCin 	DCout	6.8p
Lx	Xin	Xout	6.7p
Lin	A	2	1.22p
Lq	2	0	7.93p
Lout	q	0	31p

Kx1	Lx	L1	-0.186
Kx2	Lx	L2	-0.186
Kxd	Lx	Ld	0.190
Kd1	Ld	L1	-0.133
Kd2	Ld	L2	-0.133
Kind	Lin	Ld	5.063E-4	
Kinx	Lin	Lx	3.145E-5
Kxout	Lx	Lout	2.02E-3
Kdout	Ld	Lout	2.69E-5
Kout	Lq	Lout	0.691
.ends bfr1

.subckt branch	a	b	q
Lq	1	q	0.17p
Lb	b	1	10.4p
La	a	1	10.4p
.ends branch

.subckt split1	A	DCin	DCout	q0	q1	Xin1	Xout1
Xsplit 	splitWB	A	DCin	DCout	out	Xin1	Xout1
Xq	branch	q0	q1	out
.ends split1

VAC1	AC1	0	SIN(0 811mV 5GHz 100ps 0)
VAC2	0	AC2	SIN(0 811mV 5GHz 150ps 0)
VDC	DC1	0	PWL(0ps 0mv 20ps 1131mV)

Vin	In1	0	PWL(0ps 0mV 1ps -5mV 150ps -5mV 350ps -5mV 351ps 5mV 550ps 5mV 551ps -5mV 750ps -5mV 751ps 5mV 950ps 5mV 951ps -5mV 1150ps -5mV 1350ps -5mV 1351ps 5mV 1550ps 5mV 1750ps 5mV )

Rin	In1	1	1000	0
Rdc	DC1	d1in	1000	0	
Rx1	AC1	a1in	1000	0
Rx2	AC2	a2in	1000	0

Xsplit	split1	1	d1in	dout1	q0	q1	a1in	0
Xbfr1 	bfr1	q0	dout2	dout1	0	a2in	a2out1
Xbfr2 	bfr1	q1	0	dout2	0	a2out1 	0

.model jmod jj(rtype=1, vg=2.8mV, cap=0.064pF, r0=100, rN=17, icrit=0.1mA, Phi=pi)
.tran 0.2p 3000p 0 0.2p

.print i(Rin)
.print i(Rx1)
.print i(Rx2)
.print i(Lq|Xbfr1)
.print i(Lq|Xbfr2)

.end






