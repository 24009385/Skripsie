*KLayout buffer

.subckt	bfr1	A	dcin	dcout	q	xin	xout	
B11	4	0	jmod	area=0.5
B21	5	0	jmod	area=0.5
L1	2       4	1.98p    
L2      5	2       1.98p
Ld	DCin 	DCout	7.34p
Lx	Xin	Xout	7.28p
Lin	A	2	2.119p
Lq	2	0	7.511p
Lout	0	q	26.304p

Kx1	Lx	L1	-0.17233
Kx2	Lx	L2	-0.17233
Kxd	Lx	Ld	0.088579
Kd1	Ld	L1	-0.12779
Kd2	Ld	L2	-0.12779
Kind	Lin	Ld	2.638E-4	
Kinx	Lin	Lx	7.711E-5
Kxout	Lx	Lout	-3.194E-5
Kdout	Ld	Lout	-1.522E-5
Kout	Lq	Lout	-0.573
.ends bfr1

VAC1	AC1	0	SIN(0 811mV 5GHz 100ps 0)
VAC2	0	AC2	SIN(0 811mV 5GHz 150ps 0)
VDC	DC1	0	PWL(0ps 0mv 20ps 1131mV)

VinA	InA	0	PWL(0ps 0mV 1ps -5mV 	150ps -5mV 350ps -5mV 	351ps -5mV 550ps -5mV		551ps -5mV 750ps -5mV 		751ps -5mV 950ps -5mV 							951ps 5mV 1150ps 5mV 	1151ps 5mv 1350ps 5mV 		1351ps 5mV 1550ps 5mV 		1151ps 5mV 1750ps 5mV	1751ps -5mV)


RinA	InA	A	1000 nfree
Rdc	DC1	d1in	1000 nfree
Rx1	AC1	a1in	1000 nfree
Rx2	AC2	a2in	1000 nfree

X1	bfr1	A 	d1in	dout1	outa	a1in	a1out1
Lm1	outa	outb	1800p
X2	bfr1	outb 	dout2	dout1	out1a	a2in	a2out1
Lm2	out1a	out1b	1800p
X3	bfr1	out1b 	dout2	dout3	out2a	a1out2	a1out1
Lm3	out2a	out2b	1800p
X4	bfr1	out2b	dout4	dout3	out3a	a2out2	a2out1
Lm4	out3a	out3b	1800p
X5	bfr1	out3b	dout4	dout5	out4a	a1out2	a1out3
Lm5	out4a	out4b	1800p
X6	bfr1	out4b	dout6	dout5	out5a	a2out2	a2out3
Lm6	out5a	out5b	1800p
X7	bfr1	out5b	dout6	dout7	out6a	a1out4	a1out3
Lm7	out6a	out6b	1800p
X8	bfr1	out6b	dout8	dout7	out7	a2out4	a2out3

X9	bfr1	out7	dout8	dout9	out8	a1out4	a1out5

X10	bfr1	out8	dout10	dout9	out9	a2out4	a2out5

X11	bfr1	out9	dout10	dout11	out10	0	a1out5

X12	bfr1	out10	0	dout11	0	0	a2out5

.model jmod jj(rtype=1, vg=2.8mV, cap=0.064pF, r0=100, rN=17, icrit=0.1mA, Phi=pi)
.tran 0.2p 3000p 0 0.2p

.print i(RinA)
.print i(Lq|X2)
.print i(Lq|X3)
.print i(Lq|X4)
.print i(Lq|X5)
.print i(Lq|X6)
.print i(Lq|X7)
.print i(Lq|X8)

.end

